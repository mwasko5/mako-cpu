library ieee;
use ieee.std_logic_1164.all;

entity MEM_WB_P is
--  Port ( );
end MEM_WB_P;

architecture Behavioral of MEM_WB_P is

begin


end Behavioral;
