library ieee;
use ieee.std_logic_1164.all;

entity EX_MEM_P is
--  Port ( );
end EX_MEM_P;

architecture Behavioral of EX_MEM_P is

begin


end Behavioral;
