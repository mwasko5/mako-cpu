library ieee;
use ieee.std_logic_1164.all;

entity ID_EX_P is
--  Port ( );
end ID_EX_P;

architecture Behavioral of ID_EX_P is

begin


end Behavioral;
