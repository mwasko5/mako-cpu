library ieee;
use ieee.std_logic_1164.all;

entity IF_ID_P is
--  Port ( );
end IF_ID_P;

architecture Behavioral of IF_ID_P is

begin


end Behavioral;
